CLK = U
LED = UUUUUUUU
DIR = U
clk_div = 0000
count = 00000000
