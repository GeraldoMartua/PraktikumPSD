LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FACTORIAL IS
	PORT(	NUM	:	IN		STD_LOGIC_VECTOR(3 DOWNTO 0);
			EN		: 	IN 	STD_LOGIC;
			CLK	: 	IN		STD_LOGIC := '1';
			RES	: 	OUT 	STD_LOGIC_VECTOR(7 DOWNTO 0));
END FACTORIAL;

ARCHITECTURE MUL OF FACTORIAL IS
	SIGNAL SUM	: 	STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000001";
	SIGNAL COUNT:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";

	
	BEGIN
		PROCESS	
		BEGIN
			WAIT UNTIL CLK = '1' AND CLK'EVENT;
			IF EN = '1' THEN
				IF NUM <= "0101" THEN
					IF COUNT <= NUM THEN
						SUM <= SUM(4 DOWNTO 0)*COUNT(2 DOWNTO 0);
						COUNT <= COUNT + 1;
					END IF;
				ELSE SUM <= "00000000";
				END IF;
			END IF;
			RES <= SUM;
		END PROCESS;
		
END MUL;