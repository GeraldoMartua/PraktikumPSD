library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.Numeric_Std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ADD is
port (
	A, B		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	DATAIN		: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	ADDRESS		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLK		: IN STD_LOGIC;
	DATAOUT		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
end entity ADD;

ARCHITECTURE BEV OF ADD IS
	TYPE MEM IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL MEMORY: MEM;
	SIGNAL ADDR: INTEGER RANGE 0 TO 31;
	SIGNAL HASIL : STD_LOGIC_VECTOR(3 DOWNTO 0);
	BEGIN
	PROCESS(ADDRESS, DATAIN, CLK)
	BEGIN
		ADDR<=CONV_INTEGER(ADDRESS);
		IF (RISING_EDGE(CLK)) THEN
			HASIL <= A + B;
			DATAIN <= HASIL;
		END IF;
		MEMORY(ADDR)<=DATAIN;
		DATAOUT <= MEMORY(ADDR);
	END PROCESS;
END ARCHITECTURE BEV;