library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.Numeric_Std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity RAM_kali is
  port (
   DATAIN		: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLK			: IN STD_LOGIC;
	ADDRESS		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	W_R			: IN STD_LOGIC;
	DATA1, DATA2: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	DATAOUT		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
end entity RAM_kali;

ARCHITECTURE BEHAV OF RAM_kali IS
	TYPE MEM IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL MEMORY: MEM;
	SIGNAL ADDR: INTEGER RANGE 0 TO 31;
	SIGNAL HASIL : STD_LOGIC_VECTOR(3 DOWNTO 0);	
	BEGIN
	PROCESS(ADDRESS, DATAIN, W_R, CLK)
	BEGIN
		ADDR<=CONV_INTEGER(ADDRESS);
	IF (RISING_EDGE(CLK)) THEN	
		IF(W_R='1') THEN
			HASIL <= DATA1 * DATA2;
			DATAIN <= HASIL;
		END IF;
	END IF;
		MEMORY(ADDR)<=DATAIN;
		DATAOUT <= MEMORY(ADDR);
	END PROCESS;
END ARCHITECTURE BEHAV;