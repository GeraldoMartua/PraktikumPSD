library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.Numeric_Std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ADD is
  port (
    	MEMODATA	: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	ADDRESS		: INTEGER RANGE 0 TO 31;
	CLOCK		: IN STD_LOGIC;
	INPUT1, INPUT2	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	DATAOUT		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
end entity ADD;

ARCHITECTURE BEV OF ADD IS
	TYPE MEM IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL MEMORY: MEM;
	SIGNAL RESULT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	BEGIN
	PROCESS(ADDRESS, MEMODATA, CLOCK)
	BEGIN
		IF(CLOCK='1') THEN
			RESULT <= INPUT1 + INPUT2;
			MEMODATA <= RESULT;
			MEMORY(ADDRESS)<=MEMODATA;
		END IF;
		DATAOUT <= MEMORY(ADDRESS);
	END PROCESS;
END ARCHITECTURE BEV;