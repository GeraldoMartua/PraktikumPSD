LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY VENDINGM IS
	PORT (
	MONEY	: IN STD_LOGIC_VECTOR (2 DOWNTO 0) := "000"
	);
END VENDINGM;


ARCHITECTURE ASM OF VENDINGM IS
	TYPE S_TYPE IS (IDLE, CHECK, EJECT);
	CONSTANT COST : STD_LOGIC_VECTOR (2 DOWNTO 0) := "101";
	SIGNAL CLOCK : STD_LOGIC := '1';
	SIGNAL INPUT, SUFF, OUTPUT	: STD_LOGIC := '0';
	SIGNAL SET	: STD_LOGIC := '1';
	SIGNAL SUM, UANG : STD_LOGIC_VECTOR (2 DOWNTO 0) := "000";
	SIGNAL STATE, NSTATE	: S_TYPE;

BEGIN
	SUFF <= '0' WHEN SUM < COST ELSE
	       '1';
	INPUT <= '1' WHEN SUM > "000" ELSE
		 '0';

	PROCESS
	BEGIN
		WAIT UNTIL RISING_EDGE(CLOCK);
		IF OUTPUT = '1' THEN
			UANG <= "000";
			SUM <= SUM - COST;
		ELSE
			UANG <= MONEY;
			IF SUFF = '0' AND UANG > "000" THEN
				SUM <= SUM + UANG;
			ELSE SUM <= SUM;
			END IF;
		END IF;
		STATE <= NSTATE;
	END PROCESS;

	PROCESS (INPUT, SET, SUFF, STATE)
	BEGIN
		CASE STATE IS
		WHEN IDLE =>
			OUTPUT <= '0';
			IF INPUT = '1' THEN NSTATE <= CHECK;
			ELSE NSTATE <= IDLE;
			END IF;
		WHEN CHECK =>
			IF SET = '0' THEN NSTATE <= CHECK;
			ELSIF SUFF = '0' THEN NSTATE <= CHECK;
			ELSE NSTATE <= EJECT;
			END IF;
		WHEN EJECT =>
			NSTATE <= IDLE;
			OUTPUT <= '1';
		END CASE;
	END PROCESS;

END ASM;

	