LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CLOCK_DIVIDER IS

PORT( 	CLOCK_IN		:IN STD_LOGIC;
		CLOCK_OUT	:OUT STD_LOGIC										
	);


SIGNAL CLK			:STD_LOGIC;
SIGNAL COUNT			:STD_LOGIC_VECTOR(5 DOWNTO 0);

END CLOCK_DIVIDER;

ARCHITECTURE DIVIDE OF CLOCK_DIVIDER IS

BEGIN
	--COUNT <= "000000";
	CLOCK_OUT <= CLK;

PROCESS (CLOCK_IN)
	BEGIN
	IF (CLOCK_IN'EVENT AND CLOCK_IN = '1') THEN
	
		COUNT <= COUNT + 1;
		IF (COUNT >= 25) THEN
			COUNT <= "000000";
			CLK <= NOT(CLK);
		END IF;
	END IF;
END PROCESS;
END DIVIDE;