library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY VENDING IS
	PORT (CLK		:IN STD_LOGIC;
	      INA,INB,INC,UN	:IN STD_LOGIC := '0';
	      OUTM, OUTK, OUTU	:OUT STD_LOGIC 
	      );
END VENDING;

ARCHITECTURE MACHINE OF VENDING IS
TYPE STATE_TYPE IS (S0,S1,S2,S3,S4);		--S0=MENUNGGU INPUT DIMASUKKAN, S1=UANG YANG DIMASUKKAN KURANG MENUNGGU INPUT INA LAGI
										--S2=UANG YANG DIMASUKKAN LEBIH SEHINGGA MENGELUARKAN KEMBALIAN, S3=UANG YANG DIMASUKKAN PAS DAN MINUMAN DIKELUARKAN
										--S4=UANG YANG DIMASUKKAN TIDAK DIKENALI SEHINGGA DIKELUARKAN LAGI DARI VENDING MACHINE
SIGNAL STATE, NEXT_STATE : STATE_TYPE;
SIGNAL S, DONE : STD_LOGIC :='0'; 		--DONE=VENDING MACHINE SELESAI BEKERJA, S=MENANDAKAN NILAI UANG YANG DIMASUKKAN LEBIH BESAR DARI HARGA PADA VENDING MACHINE 
BEGIN

PROCESS
BEGIN
	WAIT UNTIL CLK='1' AND CLK'EVENT;
	STATE <= NEXT_STATE;
END PROCESS;

PROCESS (STATE,INA,INB,INC,UN,S)
BEGIN
  IF (DONE = '0') THEN
	CASE STATE IS
	WHEN S0 => 
			IF (INA ='1') THEN NEXT_STATE <= S1;
			ELSIF (INB ='1') THEN NEXT_STATE <= S3;
			ELSIF (INC ='1') THEN NEXT_STATE <= S2;
			ELSIF (UN ='1') THEN NEXT_STATE <= S4;
			ELSE NEXT_STATE <= S0;
			END IF;
	WHEN S1 =>
			IF (INA ='1') THEN NEXT_STATE <= S3;
			ELSE NEXT_STATE <= S1;
			END IF;
	WHEN S2 =>
			IF (S ='0') THEN NEXT_STATE <= S3;
			ELSE NEXT_STATE <= S2;
			END IF;
	WHEN S3 => 
			DONE <= '1';
			NEXT_STATE <= S0;
	WHEN S4 => 
			IF (S ='0') THEN NEXT_STATE <= S0;
			ELSE NEXT_STATE <= S4;
			END IF;
    	END CASE;
  ELSE NEXT_STATE <= S0;
  END IF;
END PROCESS;

PROCESS (STATE,INA,INB,INC,UN,S)
BEGIN	
	CASE STATE IS
	WHEN S0 =>  		
		IF (INB = '1') THEN OUTM <= '1';
		ELSIF (INC = '1') THEN 
			S <= '1';
			OUTK <= '1';
		ELSIF (UN = '1') THEN 
			S <= '1';
			OUTU <='1';
		ELSE 
			OUTM <= '0';
			OUTK <= '0';
			OUTU <= '0'; 
		END IF;
	WHEN S1 =>
		IF (INA = '1') THEN OUTM <= '1';
		ELSE OUTM <= '0';
		END IF;
	WHEN S2 => 
		IF (S = '1') THEN 
			OUTM <= '1';
			S <= '0';
		ELSE OUTM <= '0';
		END IF;
	WHEN S3 => DONE <= '1';
	WHEN S4 =>
		IF (S = '1') THEN 
			DONE <= '1';
			S <= '0';
		ELSE OUTM <= '0';
		END IF;	
	END CASE;
END PROCESS;

END MACHINE;