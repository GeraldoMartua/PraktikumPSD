library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.Numeric_Std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity RAM_CALC is
  port (
   DATAIN		: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLK			: IN STD_LOGIC;
	ADDRESS		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	W_R			: IN STD_LOGIC;
	MODE			: IN STD_LOGIC_VECTOR(1 DOWNTO 0); -- 00:TAMBAH ; 01:KURANG ; 10&11:KALI
	DATA1, DATA2: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	DATAOUT		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
end entity RAM_CALC;

ARCHITECTURE BEHAV OF RAM_CALC IS
	TYPE MEM IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL MEMORY: MEM;
	SIGNAL ADDR: INTEGER RANGE 0 TO 31;
	SIGNAL HASIL_TAMBAH : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL HASIL_KURANG : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL HASIL_KALI : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL ARITH_MODE : STD_LOGIC_VECTOR(1 DOWNTO 0);
	BEGIN
	PROCESS(ADDRESS, DATAIN, W_R, CLK)
	BEGIN
		ADDR<=CONV_INTEGER(ADDRESS);
	IF (RISING_EDGE(CLK)) THEN	
		IF(W_R='1') THEN
			HASIL_TAMBAH <= DATA1 + DATA2;
			HASIL_KURANG <= DATA1 - DATA2;
			HASIL_KALI <= DATA1 * DATA2;
		END IF;
	END IF;	
	END PROCESS;
	
			WITH MODE SELECT
				DATAIN <= 	HASIL_TAMBAH WHEN "00",
								HASIL_KURANG WHEN "01",
								HASIL_KALI(3 downto 0) WHEN	OTHERS;
		MEMORY(ADDR)<=DATAIN;
		DATAOUT <= MEMORY(ADDR);
		
END ARCHITECTURE BEHAV;