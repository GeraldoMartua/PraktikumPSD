LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PAYFSM IS
	PORT (
		KOIN : IN STD_LOGIC;
		CLK  : IN BIT);
END ENTITY;

ARCHITECTURE FSM OF PAYFSM IS
TYPE STATE_TYPE IS (IC, INN, W, D, WFA, ENDD, CO); --STATE TYPE
SIGNAL STATE, NEXT_STATE : STATE_TYPE;
SIGNAL TIO, SC, C, R, PA, INS, NC, DC : STD_LOGIC; --EVENT SIGNAL/OUTPUT SIGNAL SPECIFIC
SIGNAL ADC : STD_LOGIC; --INPUT SIGNAL SPECIFIC
SIGNAL X : STD_LOGIC;  --INPUT SIGNAL GENERAL
SIGNAL Z : STD_LOGIC; -- OUTPUT SIGNAL GENERAL
BEGIN
-- FLIP FLOP PROCESS
	PROCESS
	BEGIN
		WAIT UNTIL CLK ='1' AND CLK' EVENT;
		STATE <= NEXT_STATE;
	END PROCESS;

-- PAYPHONE NEXT STATE PROCESS
	PROCESS (STATE, X)
	BEGIN
	CASE STATE IS
		WHEN IC =>
			IF (X='0') THEN NEXT_STATE<=IC;
			ELSIF (X='1') THEN NEXT_STATE<=INN;
			ELSIF (ADC='1') THEN NEXT_STATE<=CO;
			ELSE NULL;
			END IF;
		WHEN INN =>
			IF (X='0') THEN NEXT_STATE <= IC;
			ELSE NEXT_STATE <= W;
			END IF;
		WHEN W => 
			IF (X='0') THEN NEXT_STATE <= IC;
			ELSE NEXT_STATE <= D;
			END IF;
		WHEN D =>
			IF (X='0') THEN NEXT_STATE <= IC;
			ELSE NEXT_STATE <= WFA;
			END IF;
		WHEN WFA =>
			IF (X='0') THEN NEXT_STATE <= IC;
			ELSE NEXT_STATE <= CO;
			END IF;
		WHEN CO =>
			IF (X='0') THEN NEXT_STATE <= IC;
			ELSE NEXT_STATE <= ENDD;
			END IF;
		WHEN ENDD =>
			NULL;
	END CASE;
END PROCESS;
-- PAYPHONE OUTPUT
	PROCESS (STATE, X)
	BEGIN
	CASE STATE IS 
		WHEN IC =>
			IF (X='0') THEN INS <= '1';
			ELSIF (X='1') THEN Z <= '0';
			ELSIF (ADC ='1') THEN NC <= '1';
			ELSE NULL;
			END IF;
		WHEN INN =>
			IF (X='0') THEN TIO <='1';
			ELSE C <= '1';
			END IF;
		WHEN W =>
			IF (X = '0') THEN TIO <='1';
			ELSE SC <= '1';
			END IF;
		WHEN D => 
			IF (X = '0') THEN TIO <='1';
			ELSE R <= '1';
			END IF;
		WHEN WFA => 
			IF (X = '0') THEN TIO <='1';
			ELSE PA <= '1';
			END IF;
		WHEN CO =>
			IF (X = '0') THEN TIO <='1';
			ELSE DC <= '1';
			END IF;
		WHEN ENDD =>
			NULL;
	END CASE;
END PROCESS;
END ARCHITECTURE;
