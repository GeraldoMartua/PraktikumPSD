LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY TELP_TB IS
END ENTITY;	

ARCHITECTURE TELP OF TELP_TB IS
SIGNAL CLK : STD_LOGIC;
SIGNAL ANGKAT : STD_LOGIC;
SIGNAL COIN : STD_LOGIC;
SIGNAL SELESAIINPUT : STD_LOGIC;
SIGNAL inputan : std_logic;
SIGNAL TELEFON : STD_LOGIC;
SIGNAL DURASI : INTEGER;
BEGIN
KONEKSI: ENTITY WORK.PUBLIC(KOIN)
PORT MAP( 	CLK=>CLK,
		ANGKAT => ANGKAT,
		COIN => COIN,
		SELESAIINPUT => SELESAIINPUT,
		INPUTAN => INPUTAN,
		TELEFON => TELEFON,
		DURASI => DURASI);

PROCESS IS
BEGIN
CLK <='1';
WAIT FOR 1 NS;
CLK <='0';
WAIT FOR 1 NS;
END PROCESS;
END ARCHITECTURE;
