LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Multiply IS
	PORT(	NUM1, NUM2	:	IN		STD_LOGIC_VECTOR(3 DOWNTO 0);
			CLK	: 	IN		STD_LOGIC := '1';
			EN		:	IN		STD_LOGIC;
			RES	: 	OUT 	STD_LOGIC_VECTOR(7 DOWNTO 0));
END Multiply;

ARCHITECTURE MULTI OF Multiply IS
	SIGNAL SUM	: 	STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
	BEGIN
		PROCESS	
		BEGIN
			WAIT UNTIL CLK = '1' AND CLK'EVENT;
			IF EN = '1' THEN
				SUM <= NUM1*NUM2;
			END IF;
		END PROCESS;
		RES <= SUM;		
END MULTI;