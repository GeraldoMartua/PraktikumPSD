LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY UpDownCounter IS
	PORT(
	RESET		: IN STD_LOGIC := '0';
	LOAD		: IN STD_LOGIC := '0';
	DIR		: IN STD_LOGIC := '0';	
	NUMBER		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	SEVSEG		: OUT STD_LOGIC_VECTOR (6 DOWNTO 0) := "0000000");
END UpDownCounter;

ARCHITECTURE Behaviour OF UpDownCounter IS
	CONSTANT CLK_FRQ	: INTEGER := 100e6;
	CONSTANT CLK_PRD	: TIME := 1000 ms / CLK_FRQ;
	SIGNAL CLK		: STD_LOGIC := '0';
	SIGNAL TEMP		: STD_LOGIC_VECTOR (3 DOWNTO 0) := "0000";

BEGIN
	CLK <= NOT CLK AFTER CLK_PRD / 2;
	
	PROCESS (CLK, RESET, LOAD, DIR, NUMBER)
	BEGIN
		IF RESET = '1'
			THEN TEMP <= "0000";
		ELSIF LOAD = '1'
			THEN TEMP <= NUMBER;
		ELSIF (RISING_EDGE(CLK))
			THEN IF TEMP = "1001"
				THEN TEMP <= "0000";
			ELSIF DIR = '0'
				THEN TEMP <= TEMP + 1;
			ELSIF DIR = '1'
				THEN TEMP <= TEMP - 1;
			END IF;
		END IF;

	END PROCESS;
	
	SEVSEG <= "1111110" WHEN TEMP = "0000" ELSE
		"0110000" WHEN TEMP = "0001" ELSE
		"1101101" WHEN TEMP = "0010" ELSE
		"1111001" WHEN TEMP = "0011" ELSE
		"0110011" WHEN TEMP = "0100" ELSE
		"1011011" WHEN TEMP = "0101" ELSE
		"0011111" WHEN TEMP = "0110" ELSE
		"1110000" WHEN TEMP = "0111" ELSE
		"1111111" WHEN TEMP = "1000" ELSE
		"1110011" WHEN TEMP = "1001";

	
END Behaviour;
